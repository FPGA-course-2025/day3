module 	notm (
		input wire A,
		output wire B
	);
 
	assign B = ~ A;

endmodule
