always  @ (a or b or sel)
begin
	... 
end
